module and_1_bit (a,b,c);

input a,b;
output c;

and and1(c,a,b);

endmodule
