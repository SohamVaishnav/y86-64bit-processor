module ALU_64_bit_tb;

reg [63:0] A,B;
wire [63:0] C,D,X,Y,Z,W,an,E,P;
wire [62:0] S;
wire SIGN,OVER;
reg S0,S1;

decoder_4_1 m1(.s0(S0),.s1(S1),.out0(E[0]),.out1(E[1]),.out2(E[2]),.out3(E[3]));

enable_64_bit i1(.e(~S0),.a(A),.b(B),.c(C),.d(D));
enable_64_bit i2(.e(E[2]),.a(A),.b(B),.c(X),.d(Y));
enable_64_bit i3(.e(E[3]),.a(A),.b(B),.c(Z),.d(W));

add_sub_64_bit a1(.a(C),.b(D),.m(S1),.sum(S),.over(OVER),.sign(SIGN));

and_64_bit f1(.a(X),.b(Y),.c(an));

xor_64_bit p1(.a(Z),.b(W),.c(P));

always@(S0,S1,A,B)
begin
    $display("S0 = %d, S1= %d, A = %b, B = %b, Sum/Difference = %b, Sign= %d, Overflow = %d, AND= %b , XOR = %b",S0,S1,A,B,S,SIGN,OVER,an,P);
end

initial
begin
    S0 = 0; S1 = 0; A = 64'b1000101111101001010110101101100101110110111110100101101101110000; B = 64'b1101110101010101100100101101110110101100110101011011100101011010;
    #10 S0 = 0; S1 = 0; A = 64'b1110011011101101101110010101110101111010101101011101110101000101; B = 64'b1011100101100010110101101010101010101110101101011101011011101110;
    #10 S0 = 0; S1 = 0; A = 64'b1100101011100101010010110101011101101101011101111111010100011011; B = 64'b1001010101110011100100101101011010101110100110101111101101100100;
    #10 S0 = 0; S1 = 1; A = 64'b1000101111101001010110101101100101110110111110100101101101110000; B = 64'b1101110101010101100100101101110110101100110101011011100101011010;
    #10 S0 = 0; S1 = 1; A = 64'b1110011011101101101110010101110101111010101101011101110101000101; B = 64'b1011100101100010110101101010101010101110101101011101011011101110;
    #10 S0 = 0; S1 = 1; A = 64'b1100101011100101010010110101011101101101011101111111010100011011; B = 64'b1001010101110011100100101101011010101110100110101111101101100100;
    #10 S0 = 1; S1 = 0; A = 64'b1000101111101001010110101101100101110110111110100101101101110000; B = 64'b1101110101010101100100101101110110101100110101011011100101011010;
    #10 S0 = 1; S1 = 0; A = 64'b1110011011101101101110010101110101111010101101011101110101000101; B = 64'b1011100101100010110101101010101010101110101101011101011011101110;
    #10 S0 = 1; S1 = 0; A = 64'b1100101011100101010010110101011101101101011101111111010100011011; B = 64'b1001010101110011100100101101011010101110100110101111101101100100;
    #10 S0 = 1; S1 = 1; A = 64'b1000101111101001010110101101100101110110111110100101101101110000; B = 64'b1101110101010101100100101101110110101100110101011011100101011010;
    #10 S0 = 1; S1 = 1; A = 64'b1110011011101101101110010101110101111010101101011101110101000101; B = 64'b1011100101100010110101101010101010101110101101011101011011101110;
    #10 S0 = 1; S1 = 1; A = 64'b1100101011100101010010110101011101101101011101111111010100011011; B = 64'b1001010101110011100100101101011010101110100110101111101101100100;
end

endmodule

