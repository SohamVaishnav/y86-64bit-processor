module enable_1_bit(e,a,out);

input e,a;
output out;

and and1(out,e,a);

endmodule


